`timescale 1ns / 1ps
// Verilog code for 16-bit single cycle MIPS CPU  
module mips_16(
    input clk,
    input reset,  
    output [15:0] pc_out,
    output [15:0] alu_result,
    output [15:0]reg3,
    output [15:0]reg4,
    output [15:0]reg5,
    output [15:0]reg2  
);  

    // Program Counter
    reg [15:0] pc_current;  
    wire signed [15:0] pc_next, pc2;  

    // Instruction
    wire [15:0] instr;  

    // Control signals
    wire [1:0] reg_dst, mem_to_reg, alu_op;  
    wire jump, branch, mem_read, mem_write, alu_src, reg_write;  
    wire sign_or_zero;

    // Register file wires
    wire [2:0] reg_write_dest;  
    wire [15:0] reg_write_data;  
    wire [2:0] reg_read_addr_1;  
    wire [15:0] reg_read_data_1;  
    wire [2:0] reg_read_addr_2;  
    wire [15:0] reg_read_data_2;  

    // ALU and immediate wires
    wire [15:0] sign_ext_im, zero_ext_im, imm_ext, read_data2;  
    wire JRControl;  
    wire [2:0] ALU_Control;  
    wire [15:0] ALU_out;  
    wire zero_flag;  
    wire signed [15:0] im_shift_1, PC_j, PC_beq, PC_4beq, PC_4beqj, PC_jr;  
    wire beq_control;  
    wire [14:0] jump_shift_1;  
    wire [15:0] mem_read_data;  
    wire [15:0] no_sign_ext;  

    // Program Counter logic
    always @(posedge clk or posedge reset) begin   
        if (reset)   
            pc_current <= 16'd0;  
        else  
            pc_current <= pc_next;  
    end  

    // PC + 2
    assign pc2 = pc_current + 16'd2;  

    // Instruction memory
    instr_mem instruction_memory(
        .pc(pc_current),
        .instruction(instr)
    );  

    // Jump shift left by 1
    assign jump_shift_1 = {instr[13:0], 1'b0};  

    // Control unit
    control control_unit(
        .reset(reset),
        .opcode(instr[15:13]),
        .reg_dst(reg_dst),
        .mem_to_reg(mem_to_reg),
        .alu_op(alu_op),
        .jump(jump),
        .branch(branch),
        .mem_read(mem_read),
        .mem_write(mem_write),
        .alu_src(alu_src),
        .reg_write(reg_write),
        .sign_or_zero(sign_or_zero)
    );  

    // Multiplexer reg_dest
    assign reg_write_dest = (reg_dst == 2'b10) ? 3'b111 : 
                            ((reg_dst == 2'b01) ? instr[6:4] : instr[9:7]);  

    // Register file
    assign reg_read_addr_1 = instr[12:10];  
    assign reg_read_addr_2 = instr[9:7];  

    register_file reg_file(
        .clk(clk),
        .rst(reset),
        .reg_write_en(reg_write),
        .reg_write_dest(reg_write_dest),
        .reg_write_data(reg_write_data),
        .reg_read_addr_1(reg_read_addr_1),
        .reg_read_data_1(reg_read_data_1),
        .reg_read_addr_2(reg_read_addr_2),
        .reg_read_data_2(reg_read_data_2),
        .reg3(reg3),
        .reg4(reg4),
        .reg5(reg5),
        .reg2(reg2)
    );  

    // Sign extend
    assign sign_ext_im = {{9{instr[6]}}, instr[6:0]};  
    assign zero_ext_im = {{9{1'b0}}, instr[6:0]};  
    assign imm_ext = (sign_or_zero == 1'b1) ? sign_ext_im : zero_ext_im;  

    // JR control
    JR_Control JRControl_unit(
        .alu_op(alu_op),
        .funct(instr[3:0]),
        .JRControl(JRControl)
    );       

    // ALU control unit
    ALUControl ALU_Control_unit(
        .ALUOp(alu_op),
        .Function(instr[3:0]),
        .ALU_Control(ALU_Control)
    );  

    // Multiplexer ALU source
    assign read_data2 = (alu_src == 1'b1) ? imm_ext : reg_read_data_2;  

    // ALU
    alu alu_unit(
        .a(reg_read_data_1),
        .b(read_data2),
        .alu_control(ALU_Control),
        .result(ALU_out),
        .zero(zero_flag)
    );  

    // Immediate shift left 1
    assign im_shift_1 = {imm_ext[14:0], 1'b0};  
    assign no_sign_ext = ~(im_shift_1) + 1'b1;  

    // PC for branch
    assign PC_beq = (im_shift_1[15] == 1'b1) ? (pc2 - no_sign_ext) : (pc2 + im_shift_1);  
    assign beq_control = branch & zero_flag;  
    assign PC_4beq = (beq_control == 1'b1) ? PC_beq : pc2;  

    // PC for jump
    assign PC_j = {pc2[15], jump_shift_1};  
    assign PC_4beqj = (jump == 1'b1) ? PC_j : PC_4beq;  
    assign PC_jr = reg_read_data_1;  

    // Next PC
    assign pc_next = (JRControl == 1'b1) ? PC_jr : PC_4beqj;  

    // Data memory
    data_memory datamem(
        .clk(clk),
        .mem_access_addr(ALU_out),
        .mem_write_data(reg_read_data_2),
        .mem_write_en(mem_write),
        .mem_read(mem_read),
        .mem_read_data(mem_read_data)
    );  

    // Write back
    assign reg_write_data = (mem_to_reg == 2'b10) ? pc2 : 
                            ((mem_to_reg == 2'b01) ? mem_read_data : ALU_out);  

    // Outputs
    assign pc_out = pc_current;  
    assign alu_result = ALU_out;  

endmodule
